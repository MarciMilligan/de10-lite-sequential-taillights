parameter IDLE      = 3'b000;
parameter HZRD      = 3'b001;
parameter SIG_L     = 3'b010;
parameter SIG_R     = 3'b011;
parameter BRK       = 3'b100;
parameter BRK_SIG_L = 3'b101;
parameter BRK_SIG_R = 3'b110;
